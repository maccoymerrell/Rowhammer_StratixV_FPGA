// asmi.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module asmi (
		input  wire [31:0] addr,          //          addr.addr
		input  wire        bulk_erase,    //    bulk_erase.bulk_erase
		output wire        busy,          //          busy.busy
		input  wire        clkin,         //         clkin.clk
		output wire        data_valid,    //    data_valid.data_valid
		input  wire [7:0]  datain,        //        datain.datain
		output wire [7:0]  dataout,       //       dataout.dataout
		input  wire        en4b_addr,     //     en4b_addr.en4b_addr
		input  wire        fast_read,     //     fast_read.fast_read
		output wire        illegal_erase, // illegal_erase.illegal_erase
		output wire        illegal_write, // illegal_write.illegal_write
		input  wire        rden,          //          rden.rden
		output wire [7:0]  rdid_out,      //      rdid_out.rdid_out
		input  wire        read_rdid,     //     read_rdid.read_rdid
		input  wire        read_status,   //   read_status.read_status
		input  wire        reset,         //         reset.reset
		input  wire        shift_bytes,   //   shift_bytes.shift_bytes
		output wire [7:0]  status_out,    //    status_out.status_out
		input  wire        wren,          //          wren.wren
		input  wire        write          //         write.write
	);

	asmi_asmi_parallel_0 asmi_parallel_0 (
		.clkin         (clkin),         //         clkin.clk
		.fast_read     (fast_read),     //     fast_read.fast_read
		.rden          (rden),          //          rden.rden
		.addr          (addr),          //          addr.addr
		.read_status   (read_status),   //   read_status.read_status
		.write         (write),         //         write.write
		.datain        (datain),        //        datain.datain
		.shift_bytes   (shift_bytes),   //   shift_bytes.shift_bytes
		.bulk_erase    (bulk_erase),    //    bulk_erase.bulk_erase
		.wren          (wren),          //          wren.wren
		.read_rdid     (read_rdid),     //     read_rdid.read_rdid
		.en4b_addr     (en4b_addr),     //     en4b_addr.en4b_addr
		.reset         (reset),         //         reset.reset
		.dataout       (dataout),       //       dataout.dataout
		.busy          (busy),          //          busy.busy
		.data_valid    (data_valid),    //    data_valid.data_valid
		.status_out    (status_out),    //    status_out.status_out
		.illegal_write (illegal_write), // illegal_write.illegal_write
		.illegal_erase (illegal_erase), // illegal_erase.illegal_erase
		.rdid_out      (rdid_out)       //      rdid_out.rdid_out
	);

endmodule
