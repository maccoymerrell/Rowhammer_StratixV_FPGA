// pcie_hip_avmm.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module pcie_hip_avmm (
		output wire [7:0]   avl_to_asmi_0_conduit_end_sfl_address,       // avl_to_asmi_0_conduit_end.sfl_address
		output wire         avl_to_asmi_0_conduit_end_sfl_read,          //                          .sfl_read
		input  wire [31:0]  avl_to_asmi_0_conduit_end_sfl_readdata_from, //                          .sfl_readdata_from
		output wire         avl_to_asmi_0_conduit_end_sfl_write,         //                          .sfl_write
		output wire [31:0]  avl_to_asmi_0_conduit_end_sfl_writedata_to,  //                          .sfl_writedata_to
		output wire         avl_to_asmi_0_conduit_end_sfl_clk,           //                          .sfl_clk
		output wire         avl_to_asmi_0_conduit_end_sfl_reset,         //                          .sfl_reset
		input  wire         clk_clk,                                     //                       clk.clk
		input  wire         clk_1_clk,                                   //                     clk_1.clk
		input  wire [31:0]  fast_mem_address,                            //                  fast_mem.address
		input  wire         fast_mem_read,                               //                          .read
		output wire [511:0] fast_mem_readdata,                           //                          .readdata
		output wire         fast_mem_readdatavalid,                      //                          .readdatavalid
		output wire         fast_mem_waitrequest,                        //                          .waitrequest
		input  wire         fast_mem_write,                              //                          .write
		input  wire [511:0] fast_mem_writedata,                          //                          .writedata
		input  wire [5:0]   fast_mem_burstcount,                         //                          .burstcount
		input  wire         fast_mem_lock,                               //                          .lock
		input  wire [31:0]  hip_ctrl_test_in,                            //                  hip_ctrl.test_in
		input  wire         hip_ctrl_simu_mode_pipe,                     //                          .simu_mode_pipe
		input  wire         hip_serial_rx_in0,                           //                hip_serial.rx_in0
		input  wire         hip_serial_rx_in1,                           //                          .rx_in1
		input  wire         hip_serial_rx_in2,                           //                          .rx_in2
		input  wire         hip_serial_rx_in3,                           //                          .rx_in3
		output wire         hip_serial_tx_out0,                          //                          .tx_out0
		output wire         hip_serial_tx_out1,                          //                          .tx_out1
		output wire         hip_serial_tx_out2,                          //                          .tx_out2
		output wire         hip_serial_tx_out3,                          //                          .tx_out3
		output wire [12:0]  memory_mem_a,                                //                    memory.mem_a
		output wire [2:0]   memory_mem_ba,                               //                          .mem_ba
		output wire [1:0]   memory_mem_ck,                               //                          .mem_ck
		output wire [1:0]   memory_mem_ck_n,                             //                          .mem_ck_n
		output wire [1:0]   memory_mem_cke,                              //                          .mem_cke
		output wire [1:0]   memory_mem_cs_n,                             //                          .mem_cs_n
		output wire [7:0]   memory_mem_dm,                               //                          .mem_dm
		output wire [0:0]   memory_mem_ras_n,                            //                          .mem_ras_n
		output wire [0:0]   memory_mem_cas_n,                            //                          .mem_cas_n
		output wire [0:0]   memory_mem_we_n,                             //                          .mem_we_n
		output wire         memory_mem_reset_n,                          //                          .mem_reset_n
		inout  wire [63:0]  memory_mem_dq,                               //                          .mem_dq
		inout  wire [7:0]   memory_mem_dqs,                              //                          .mem_dqs
		inout  wire [7:0]   memory_mem_dqs_n,                            //                          .mem_dqs_n
		output wire [1:0]   memory_mem_odt,                              //                          .mem_odt
		output wire [12:0]  memory_1_mem_a,                              //                  memory_1.mem_a
		output wire [2:0]   memory_1_mem_ba,                             //                          .mem_ba
		output wire [1:0]   memory_1_mem_ck,                             //                          .mem_ck
		output wire [1:0]   memory_1_mem_ck_n,                           //                          .mem_ck_n
		output wire [1:0]   memory_1_mem_cke,                            //                          .mem_cke
		output wire [1:0]   memory_1_mem_cs_n,                           //                          .mem_cs_n
		output wire [7:0]   memory_1_mem_dm,                             //                          .mem_dm
		output wire [0:0]   memory_1_mem_ras_n,                          //                          .mem_ras_n
		output wire [0:0]   memory_1_mem_cas_n,                          //                          .mem_cas_n
		output wire [0:0]   memory_1_mem_we_n,                           //                          .mem_we_n
		output wire         memory_1_mem_reset_n,                        //                          .mem_reset_n
		inout  wire [63:0]  memory_1_mem_dq,                             //                          .mem_dq
		inout  wire [7:0]   memory_1_mem_dqs,                            //                          .mem_dqs
		inout  wire [7:0]   memory_1_mem_dqs_n,                          //                          .mem_dqs_n
		output wire [1:0]   memory_1_mem_odt,                            //                          .mem_odt
		input  wire         mgmt_clk_clk,                                //                  mgmt_clk.clk
		input  wire         mgmt_rst_reset,                              //                  mgmt_rst.reset
		input  wire         oct_rzqin,                                   //                       oct.rzqin
		input  wire         oct_1_rzqin,                                 //                     oct_1.rzqin
		input  wire         pcie_npor_npor,                              //                 pcie_npor.npor
		input  wire         pcie_npor_pin_perst,                         //                          .pin_perst
		input  wire         pcie_refclock_clk,                           //             pcie_refclock.clk
		input  wire         reconfig_xcvr_clk_clk,                       //         reconfig_xcvr_clk.clk
		input  wire         reconfig_xcvr_rst_reset,                     //         reconfig_xcvr_rst.reset
		input  wire         reset_reset_n,                               //                     reset.reset_n
		input  wire         reset_1_reset_n,                             //                   reset_1.reset_n
		input  wire [31:0]  slow_mem_address,                            //                  slow_mem.address
		input  wire         slow_mem_read,                               //                          .read
		output wire [511:0] slow_mem_readdata,                           //                          .readdata
		output wire         slow_mem_readdatavalid,                      //                          .readdatavalid
		input  wire         slow_mem_write,                              //                          .write
		input  wire [511:0] slow_mem_writedata,                          //                          .writedata
		output wire         slow_mem_waitrequest,                        //                          .waitrequest
		input  wire [5:0]   slow_mem_burstcount,                         //                          .burstcount
		input  wire         slow_mem_lock                                //                          .lock
	);

	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_readdata;               // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> pcie_reconfig_driver_0:reconfig_mgmt_readdata
	wire          pcie_reconfig_driver_0_reconfig_mgmt_waitrequest;            // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> pcie_reconfig_driver_0:reconfig_mgmt_waitrequest
	wire    [6:0] pcie_reconfig_driver_0_reconfig_mgmt_address;                // pcie_reconfig_driver_0:reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          pcie_reconfig_driver_0_reconfig_mgmt_read;                   // pcie_reconfig_driver_0:reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire          pcie_reconfig_driver_0_reconfig_mgmt_write;                  // pcie_reconfig_driver_0:reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_writedata;              // pcie_reconfig_driver_0:reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire          dut_coreclkout_clk;                                          // DUT:coreclkout -> [avl_to_asmi_0:clk, irq_mapper:clk, mm_interconnect_0:DUT_coreclkout_clk, mm_interconnect_1:DUT_coreclkout_clk, mm_interconnect_2:DUT_coreclkout_clk, pcie_reconfig_driver_0:pld_clk, rst_controller:clk]
	wire    [1:0] dut_hip_currentspeed_currentspeed;                           // DUT:currentspeed -> pcie_reconfig_driver_0:currentspeed
	wire          dut_hip_status_derr_cor_ext_rcv;                             // DUT:derr_cor_ext_rcv -> pcie_reconfig_driver_0:derr_cor_ext_rcv_drv
	wire          dut_hip_status_hotrst_exit;                                  // DUT:hotrst_exit -> pcie_reconfig_driver_0:hotrst_exit_drv
	wire          dut_hip_status_rx_par_err;                                   // DUT:rx_par_err -> pcie_reconfig_driver_0:rx_par_err_drv
	wire   [11:0] dut_hip_status_ko_cpl_spc_data;                              // DUT:ko_cpl_spc_data -> pcie_reconfig_driver_0:ko_cpl_spc_data_drv
	wire          dut_hip_status_dlup_exit;                                    // DUT:dlup_exit -> pcie_reconfig_driver_0:dlup_exit_drv
	wire          dut_hip_status_derr_cor_ext_rpl;                             // DUT:derr_cor_ext_rpl -> pcie_reconfig_driver_0:derr_cor_ext_rpl_drv
	wire          dut_hip_status_l2_exit;                                      // DUT:l2_exit -> pcie_reconfig_driver_0:l2_exit_drv
	wire          dut_hip_status_dlup;                                         // DUT:dlup -> pcie_reconfig_driver_0:dlup_drv
	wire    [3:0] dut_hip_status_int_status;                                   // DUT:int_status -> pcie_reconfig_driver_0:int_status_drv
	wire          dut_hip_status_ev128ns;                                      // DUT:ev128ns -> pcie_reconfig_driver_0:ev128ns_drv
	wire    [4:0] dut_hip_status_ltssmstate;                                   // DUT:ltssmstate -> pcie_reconfig_driver_0:ltssmstate_drv
	wire    [1:0] dut_hip_status_tx_par_err;                                   // DUT:tx_par_err -> pcie_reconfig_driver_0:tx_par_err_drv
	wire    [3:0] dut_hip_status_lane_act;                                     // DUT:lane_act -> pcie_reconfig_driver_0:lane_act_drv
	wire          dut_hip_status_cfg_par_err;                                  // DUT:cfg_par_err -> pcie_reconfig_driver_0:cfg_par_err_drv
	wire          dut_hip_status_derr_rpl;                                     // DUT:derr_rpl -> pcie_reconfig_driver_0:derr_rpl_drv
	wire          dut_hip_status_ev1us;                                        // DUT:ev1us -> pcie_reconfig_driver_0:ev1us_drv
	wire    [7:0] dut_hip_status_ko_cpl_spc_header;                            // DUT:ko_cpl_spc_header -> pcie_reconfig_driver_0:ko_cpl_spc_header_drv
	wire          alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy;             // alt_xcvr_reconfig_0:reconfig_busy -> pcie_reconfig_driver_0:reconfig_busy
	wire  [275:0] dut_reconfig_from_xcvr_reconfig_from_xcvr;                   // DUT:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [419:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr;       // alt_xcvr_reconfig_0:reconfig_to_xcvr -> DUT:reconfig_to_xcvr
	wire          dut_rxm_bar0_waitrequest;                                    // mm_interconnect_0:DUT_Rxm_BAR0_waitrequest -> DUT:RxmWaitRequest_0_i
	wire  [127:0] dut_rxm_bar0_readdata;                                       // mm_interconnect_0:DUT_Rxm_BAR0_readdata -> DUT:RxmReadData_0_i
	wire   [63:0] dut_rxm_bar0_address;                                        // DUT:RxmAddress_0_o -> mm_interconnect_0:DUT_Rxm_BAR0_address
	wire          dut_rxm_bar0_read;                                           // DUT:RxmRead_0_o -> mm_interconnect_0:DUT_Rxm_BAR0_read
	wire   [15:0] dut_rxm_bar0_byteenable;                                     // DUT:RxmByteEnable_0_o -> mm_interconnect_0:DUT_Rxm_BAR0_byteenable
	wire          dut_rxm_bar0_readdatavalid;                                  // mm_interconnect_0:DUT_Rxm_BAR0_readdatavalid -> DUT:RxmReadDataValid_0_i
	wire          dut_rxm_bar0_write;                                          // DUT:RxmWrite_0_o -> mm_interconnect_0:DUT_Rxm_BAR0_write
	wire  [127:0] dut_rxm_bar0_writedata;                                      // DUT:RxmWriteData_0_o -> mm_interconnect_0:DUT_Rxm_BAR0_writedata
	wire    [5:0] dut_rxm_bar0_burstcount;                                     // DUT:RxmBurstCount_0_o -> mm_interconnect_0:DUT_Rxm_BAR0_burstcount
	wire          mm_interconnect_0_dut_cra_chipselect;                        // mm_interconnect_0:DUT_Cra_chipselect -> DUT:CraChipSelect_i
	wire   [31:0] mm_interconnect_0_dut_cra_readdata;                          // DUT:CraReadData_o -> mm_interconnect_0:DUT_Cra_readdata
	wire          mm_interconnect_0_dut_cra_waitrequest;                       // DUT:CraWaitRequest_o -> mm_interconnect_0:DUT_Cra_waitrequest
	wire   [13:0] mm_interconnect_0_dut_cra_address;                           // mm_interconnect_0:DUT_Cra_address -> DUT:CraAddress_i
	wire          mm_interconnect_0_dut_cra_read;                              // mm_interconnect_0:DUT_Cra_read -> DUT:CraRead
	wire    [3:0] mm_interconnect_0_dut_cra_byteenable;                        // mm_interconnect_0:DUT_Cra_byteenable -> DUT:CraByteEnable_i
	wire          mm_interconnect_0_dut_cra_write;                             // mm_interconnect_0:DUT_Cra_write -> DUT:CraWrite
	wire   [31:0] mm_interconnect_0_dut_cra_writedata;                         // mm_interconnect_0:DUT_Cra_writedata -> DUT:CraWriteData_i
	wire   [31:0] mm_interconnect_0_mem_if_ddr3_emif_1_csr_readdata;           // mem_if_ddr3_emif_1:csr_rdata -> mm_interconnect_0:mem_if_ddr3_emif_1_csr_readdata
	wire          mm_interconnect_0_mem_if_ddr3_emif_1_csr_waitrequest;        // mem_if_ddr3_emif_1:csr_waitrequest -> mm_interconnect_0:mem_if_ddr3_emif_1_csr_waitrequest
	wire   [15:0] mm_interconnect_0_mem_if_ddr3_emif_1_csr_address;            // mm_interconnect_0:mem_if_ddr3_emif_1_csr_address -> mem_if_ddr3_emif_1:csr_addr
	wire          mm_interconnect_0_mem_if_ddr3_emif_1_csr_read;               // mm_interconnect_0:mem_if_ddr3_emif_1_csr_read -> mem_if_ddr3_emif_1:csr_read_req
	wire    [3:0] mm_interconnect_0_mem_if_ddr3_emif_1_csr_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_1_csr_byteenable -> mem_if_ddr3_emif_1:csr_be
	wire          mm_interconnect_0_mem_if_ddr3_emif_1_csr_readdatavalid;      // mem_if_ddr3_emif_1:csr_rdata_valid -> mm_interconnect_0:mem_if_ddr3_emif_1_csr_readdatavalid
	wire          mm_interconnect_0_mem_if_ddr3_emif_1_csr_write;              // mm_interconnect_0:mem_if_ddr3_emif_1_csr_write -> mem_if_ddr3_emif_1:csr_write_req
	wire   [31:0] mm_interconnect_0_mem_if_ddr3_emif_1_csr_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_1_csr_writedata -> mem_if_ddr3_emif_1:csr_wdata
	wire          mem_if_ddr3_emif_1_afi_clk_clk;                              // mem_if_ddr3_emif_1:afi_clk -> [mm_interconnect_0:mem_if_ddr3_emif_1_afi_clk_clk, mm_interconnect_2:mem_if_ddr3_emif_1_afi_clk_clk, rst_controller_002:clk]
	wire   [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_csr_readdata;           // mem_if_ddr3_emif_0:csr_rdata -> mm_interconnect_0:mem_if_ddr3_emif_0_csr_readdata
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_csr_waitrequest;        // mem_if_ddr3_emif_0:csr_waitrequest -> mm_interconnect_0:mem_if_ddr3_emif_0_csr_waitrequest
	wire   [15:0] mm_interconnect_0_mem_if_ddr3_emif_0_csr_address;            // mm_interconnect_0:mem_if_ddr3_emif_0_csr_address -> mem_if_ddr3_emif_0:csr_addr
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_csr_read;               // mm_interconnect_0:mem_if_ddr3_emif_0_csr_read -> mem_if_ddr3_emif_0:csr_read_req
	wire    [3:0] mm_interconnect_0_mem_if_ddr3_emif_0_csr_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_0_csr_byteenable -> mem_if_ddr3_emif_0:csr_be
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_csr_readdatavalid;      // mem_if_ddr3_emif_0:csr_rdata_valid -> mm_interconnect_0:mem_if_ddr3_emif_0_csr_readdatavalid
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_csr_write;              // mm_interconnect_0:mem_if_ddr3_emif_0_csr_write -> mem_if_ddr3_emif_0:csr_write_req
	wire   [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_csr_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_0_csr_writedata -> mem_if_ddr3_emif_0:csr_wdata
	wire          mem_if_ddr3_emif_0_afi_clk_clk;                              // mem_if_ddr3_emif_0:afi_clk -> [mm_interconnect_0:mem_if_ddr3_emif_0_afi_clk_clk, mm_interconnect_1:mem_if_ddr3_emif_0_afi_clk_clk, rst_controller_001:clk]
	wire   [31:0] mm_interconnect_0_avl_to_asmi_0_s0_readdata;                 // avl_to_asmi_0:avs_s0_readdata -> mm_interconnect_0:avl_to_asmi_0_s0_readdata
	wire    [7:0] mm_interconnect_0_avl_to_asmi_0_s0_address;                  // mm_interconnect_0:avl_to_asmi_0_s0_address -> avl_to_asmi_0:avs_s0_address
	wire          mm_interconnect_0_avl_to_asmi_0_s0_read;                     // mm_interconnect_0:avl_to_asmi_0_s0_read -> avl_to_asmi_0:avs_s0_read
	wire          mm_interconnect_0_avl_to_asmi_0_s0_write;                    // mm_interconnect_0:avl_to_asmi_0_s0_write -> avl_to_asmi_0:avs_s0_write
	wire   [31:0] mm_interconnect_0_avl_to_asmi_0_s0_writedata;                // mm_interconnect_0:avl_to_asmi_0_s0_writedata -> avl_to_asmi_0:avs_s0_writedata
	wire          dut_rxm_bar2_waitrequest;                                    // mm_interconnect_1:DUT_Rxm_BAR2_waitrequest -> DUT:RxmWaitRequest_2_i
	wire  [127:0] dut_rxm_bar2_readdata;                                       // mm_interconnect_1:DUT_Rxm_BAR2_readdata -> DUT:RxmReadData_2_i
	wire   [63:0] dut_rxm_bar2_address;                                        // DUT:RxmAddress_2_o -> mm_interconnect_1:DUT_Rxm_BAR2_address
	wire          dut_rxm_bar2_read;                                           // DUT:RxmRead_2_o -> mm_interconnect_1:DUT_Rxm_BAR2_read
	wire   [15:0] dut_rxm_bar2_byteenable;                                     // DUT:RxmByteEnable_2_o -> mm_interconnect_1:DUT_Rxm_BAR2_byteenable
	wire          dut_rxm_bar2_readdatavalid;                                  // mm_interconnect_1:DUT_Rxm_BAR2_readdatavalid -> DUT:RxmReadDataValid_2_i
	wire          dut_rxm_bar2_write;                                          // DUT:RxmWrite_2_o -> mm_interconnect_1:DUT_Rxm_BAR2_write
	wire  [127:0] dut_rxm_bar2_writedata;                                      // DUT:RxmWriteData_2_o -> mm_interconnect_1:DUT_Rxm_BAR2_writedata
	wire    [5:0] dut_rxm_bar2_burstcount;                                     // DUT:RxmBurstCount_2_o -> mm_interconnect_1:DUT_Rxm_BAR2_burstcount
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_beginbursttransfer; // mm_interconnect_1:mem_if_ddr3_emif_0_avl_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin
	wire  [511:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_readdata;           // mem_if_ddr3_emif_0:avl_rdata -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_readdata
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_waitrequest;        // mem_if_ddr3_emif_0:avl_ready -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_waitrequest
	wire   [23:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_address;            // mm_interconnect_1:mem_if_ddr3_emif_0_avl_address -> mem_if_ddr3_emif_0:avl_addr
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_read;               // mm_interconnect_1:mem_if_ddr3_emif_0_avl_read -> mem_if_ddr3_emif_0:avl_read_req
	wire   [63:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_byteenable;         // mm_interconnect_1:mem_if_ddr3_emif_0_avl_byteenable -> mem_if_ddr3_emif_0:avl_be
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_readdatavalid;      // mem_if_ddr3_emif_0:avl_rdata_valid -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_readdatavalid
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_write;              // mm_interconnect_1:mem_if_ddr3_emif_0_avl_write -> mem_if_ddr3_emif_0:avl_write_req
	wire  [511:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_writedata;          // mm_interconnect_1:mem_if_ddr3_emif_0_avl_writedata -> mem_if_ddr3_emif_0:avl_wdata
	wire    [2:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_burstcount;         // mm_interconnect_1:mem_if_ddr3_emif_0_avl_burstcount -> mem_if_ddr3_emif_0:avl_size
	wire          dut_rxm_bar4_waitrequest;                                    // mm_interconnect_2:DUT_Rxm_BAR4_waitrequest -> DUT:RxmWaitRequest_4_i
	wire  [127:0] dut_rxm_bar4_readdata;                                       // mm_interconnect_2:DUT_Rxm_BAR4_readdata -> DUT:RxmReadData_4_i
	wire   [63:0] dut_rxm_bar4_address;                                        // DUT:RxmAddress_4_o -> mm_interconnect_2:DUT_Rxm_BAR4_address
	wire          dut_rxm_bar4_read;                                           // DUT:RxmRead_4_o -> mm_interconnect_2:DUT_Rxm_BAR4_read
	wire   [15:0] dut_rxm_bar4_byteenable;                                     // DUT:RxmByteEnable_4_o -> mm_interconnect_2:DUT_Rxm_BAR4_byteenable
	wire          dut_rxm_bar4_readdatavalid;                                  // mm_interconnect_2:DUT_Rxm_BAR4_readdatavalid -> DUT:RxmReadDataValid_4_i
	wire          dut_rxm_bar4_write;                                          // DUT:RxmWrite_4_o -> mm_interconnect_2:DUT_Rxm_BAR4_write
	wire  [127:0] dut_rxm_bar4_writedata;                                      // DUT:RxmWriteData_4_o -> mm_interconnect_2:DUT_Rxm_BAR4_writedata
	wire    [5:0] dut_rxm_bar4_burstcount;                                     // DUT:RxmBurstCount_4_o -> mm_interconnect_2:DUT_Rxm_BAR4_burstcount
	wire          mm_interconnect_2_mem_if_ddr3_emif_1_avl_beginbursttransfer; // mm_interconnect_2:mem_if_ddr3_emif_1_avl_beginbursttransfer -> mem_if_ddr3_emif_1:avl_burstbegin
	wire  [511:0] mm_interconnect_2_mem_if_ddr3_emif_1_avl_readdata;           // mem_if_ddr3_emif_1:avl_rdata -> mm_interconnect_2:mem_if_ddr3_emif_1_avl_readdata
	wire          mm_interconnect_2_mem_if_ddr3_emif_1_avl_waitrequest;        // mem_if_ddr3_emif_1:avl_ready -> mm_interconnect_2:mem_if_ddr3_emif_1_avl_waitrequest
	wire   [23:0] mm_interconnect_2_mem_if_ddr3_emif_1_avl_address;            // mm_interconnect_2:mem_if_ddr3_emif_1_avl_address -> mem_if_ddr3_emif_1:avl_addr
	wire          mm_interconnect_2_mem_if_ddr3_emif_1_avl_read;               // mm_interconnect_2:mem_if_ddr3_emif_1_avl_read -> mem_if_ddr3_emif_1:avl_read_req
	wire   [63:0] mm_interconnect_2_mem_if_ddr3_emif_1_avl_byteenable;         // mm_interconnect_2:mem_if_ddr3_emif_1_avl_byteenable -> mem_if_ddr3_emif_1:avl_be
	wire          mm_interconnect_2_mem_if_ddr3_emif_1_avl_readdatavalid;      // mem_if_ddr3_emif_1:avl_rdata_valid -> mm_interconnect_2:mem_if_ddr3_emif_1_avl_readdatavalid
	wire          mm_interconnect_2_mem_if_ddr3_emif_1_avl_write;              // mm_interconnect_2:mem_if_ddr3_emif_1_avl_write -> mem_if_ddr3_emif_1:avl_write_req
	wire  [511:0] mm_interconnect_2_mem_if_ddr3_emif_1_avl_writedata;          // mm_interconnect_2:mem_if_ddr3_emif_1_avl_writedata -> mem_if_ddr3_emif_1:avl_wdata
	wire    [2:0] mm_interconnect_2_mem_if_ddr3_emif_1_avl_burstcount;         // mm_interconnect_2:mem_if_ddr3_emif_1_avl_burstcount -> mem_if_ddr3_emif_1:avl_size
	wire   [15:0] dut_rxmirq_irq;                                              // irq_mapper:sender_irq -> DUT:RxmIrq_i
	wire          rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [avl_to_asmi_0:reset, irq_mapper:reset, mm_interconnect_0:avl_to_asmi_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:move_engine_0_rst_reset_bridge_in_reset_reset, mm_interconnect_2:move_engine_0_rst_reset_bridge_in_reset_reset]
	wire          dut_nreset_status_reset;                                     // DUT:reset_status -> rst_controller:reset_in0
	wire          rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:mem_if_ddr3_emif_0_csr_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_interconnect_0:mem_if_ddr3_emif_1_csr_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_1_soft_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mem_if_ddr3_emif_1_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mem_if_ddr3_emif_1_soft_reset_reset_bridge_in_reset_reset]

	altpcie_sv_hip_avmm_hwtcl #(
		.lane_mask_hwtcl                          ("x4"),
		.gen123_lane_rate_mode_hwtcl              ("Gen3 (8.0 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("3.0"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.in_cvp_mode_hwtcl                        (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.enable_power_on_rst_pulse_hwtcl          (0),
		.enable_pcisigtest_hwtcl                  (0),
		.bar0_size_mask_hwtcl                     (20),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Disabled"),
		.bar0_prefetchable_hwtcl                  ("Disabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (30),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Enabled"),
		.bar2_prefetchable_hwtcl                  ("Enabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (30),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Enabled"),
		.bar4_prefetchable_hwtcl                  ("Enabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (6487),
		.device_id_hwtcl                          (2387),
		.revision_id_hwtcl                        (179),
		.class_code_hwtcl                         (360448),
		.subsystem_vendor_id_hwtcl                (4277),
		.subsystem_device_id_hwtcl                (36948),
		.max_payload_size_hwtcl                   (256),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("NONE"),
		.enable_completion_timeout_disable_hwtcl  (0),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (4466),
		.vsec_rev_hwtcl                           (0),
		.user_id_hwtcl                            (0),
		.avmm_width_hwtcl                         (128),
		.AVALON_ADDR_WIDTH                        (64),
		.avmm_burst_width_hwtcl                   (6),
		.CB_PCIE_MODE                             (0),
		.CB_PCIE_RX_LITE                          (0),
		.CB_RXM_DATA_WIDTH                        (128),
		.CG_AVALON_S_ADDR_WIDTH                   (64),
		.CG_IMPL_CRA_AV_SLAVE_PORT                (1),
		.CG_ENABLE_ADVANCED_INTERRUPT             (1),
		.CG_ENABLE_A2P_INTERRUPT                  (0),
		.CB_A2P_ADDR_MAP_IS_FIXED                 (0),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES              (2),
		.BYPASSS_A2P_TRANSLATION                  (0),
		.a2p_pass_thru_bits                       (8),
		.ast_width_hwtcl                          ("Avalon-ST 128-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (248500),
		.port_width_be_hwtcl                      (16),
		.port_width_data_hwtcl                    (128),
		.hip_reconfig_hwtcl                       (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("true"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (50),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (358),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (56),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (112),
		.cpl_spc_data_hwtcl                       (448),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (420),
		.reconfig_from_xcvr_width                 (276),
		.single_rx_detect_hwtcl                   (4),
		.hip_hard_reset_hwtcl                     (0),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15)
	) dut (
		.coreclkout           (dut_coreclkout_clk),                                    //          coreclkout.clk
		.refclk               (pcie_refclock_clk),                                     //              refclk.clk
		.npor                 (pcie_npor_npor),                                        //                npor.npor
		.pin_perst            (pcie_npor_pin_perst),                                   //                    .pin_perst
		.reset_status         (dut_nreset_status_reset),                               //       nreset_status.reset_n
		.RxmAddress_0_o       (dut_rxm_bar0_address),                                  //            Rxm_BAR0.address
		.RxmRead_0_o          (dut_rxm_bar0_read),                                     //                    .read
		.RxmWaitRequest_0_i   (dut_rxm_bar0_waitrequest),                              //                    .waitrequest
		.RxmWrite_0_o         (dut_rxm_bar0_write),                                    //                    .write
		.RxmReadDataValid_0_i (dut_rxm_bar0_readdatavalid),                            //                    .readdatavalid
		.RxmReadData_0_i      (dut_rxm_bar0_readdata),                                 //                    .readdata
		.RxmWriteData_0_o     (dut_rxm_bar0_writedata),                                //                    .writedata
		.RxmBurstCount_0_o    (dut_rxm_bar0_burstcount),                               //                    .burstcount
		.RxmByteEnable_0_o    (dut_rxm_bar0_byteenable),                               //                    .byteenable
		.RxmAddress_1_o       (),                                                      //            Rxm_BAR1.address
		.RxmRead_1_o          (),                                                      //                    .read
		.RxmWaitRequest_1_i   (),                                                      //                    .waitrequest
		.RxmWrite_1_o         (),                                                      //                    .write
		.RxmReadDataValid_1_i (),                                                      //                    .readdatavalid
		.RxmReadData_1_i      (),                                                      //                    .readdata
		.RxmWriteData_1_o     (),                                                      //                    .writedata
		.RxmBurstCount_1_o    (),                                                      //                    .burstcount
		.RxmByteEnable_1_o    (),                                                      //                    .byteenable
		.RxmAddress_2_o       (dut_rxm_bar2_address),                                  //            Rxm_BAR2.address
		.RxmRead_2_o          (dut_rxm_bar2_read),                                     //                    .read
		.RxmWaitRequest_2_i   (dut_rxm_bar2_waitrequest),                              //                    .waitrequest
		.RxmWrite_2_o         (dut_rxm_bar2_write),                                    //                    .write
		.RxmReadDataValid_2_i (dut_rxm_bar2_readdatavalid),                            //                    .readdatavalid
		.RxmReadData_2_i      (dut_rxm_bar2_readdata),                                 //                    .readdata
		.RxmWriteData_2_o     (dut_rxm_bar2_writedata),                                //                    .writedata
		.RxmBurstCount_2_o    (dut_rxm_bar2_burstcount),                               //                    .burstcount
		.RxmByteEnable_2_o    (dut_rxm_bar2_byteenable),                               //                    .byteenable
		.RxmAddress_4_o       (dut_rxm_bar4_address),                                  //            Rxm_BAR4.address
		.RxmRead_4_o          (dut_rxm_bar4_read),                                     //                    .read
		.RxmWaitRequest_4_i   (dut_rxm_bar4_waitrequest),                              //                    .waitrequest
		.RxmWrite_4_o         (dut_rxm_bar4_write),                                    //                    .write
		.RxmReadDataValid_4_i (dut_rxm_bar4_readdatavalid),                            //                    .readdatavalid
		.RxmReadData_4_i      (dut_rxm_bar4_readdata),                                 //                    .readdata
		.RxmWriteData_4_o     (dut_rxm_bar4_writedata),                                //                    .writedata
		.RxmBurstCount_4_o    (dut_rxm_bar4_burstcount),                               //                    .burstcount
		.RxmByteEnable_4_o    (dut_rxm_bar4_byteenable),                               //                    .byteenable
		.RxmIrq_i             (dut_rxmirq_irq),                                        //              RxmIrq.irq
		.MsiIntfc_o           (),                                                      //       MSI_Interface.msi_intfc
		.MsiControl_o         (),                                                      //         MSI_Control.msi_control
		.MsixIntfc_o          (),                                                      //      MSIX_Interface.msix_intfc
		.IntxReq_i            (),                                                      //      INTX_Interface.intx_req
		.IntxAck_o            (),                                                      //                    .intx_ack
		.derr_cor_ext_rcv     (dut_hip_status_derr_cor_ext_rcv),                       //          hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (dut_hip_status_derr_cor_ext_rpl),                       //                    .derr_cor_ext_rpl
		.derr_rpl             (dut_hip_status_derr_rpl),                               //                    .derr_rpl
		.dlup                 (dut_hip_status_dlup),                                   //                    .dlup
		.dlup_exit            (dut_hip_status_dlup_exit),                              //                    .dlup_exit
		.ev128ns              (dut_hip_status_ev128ns),                                //                    .ev128ns
		.ev1us                (dut_hip_status_ev1us),                                  //                    .ev1us
		.hotrst_exit          (dut_hip_status_hotrst_exit),                            //                    .hotrst_exit
		.int_status           (dut_hip_status_int_status),                             //                    .int_status
		.l2_exit              (dut_hip_status_l2_exit),                                //                    .l2_exit
		.lane_act             (dut_hip_status_lane_act),                               //                    .lane_act
		.ltssmstate           (dut_hip_status_ltssmstate),                             //                    .ltssmstate
		.rx_par_err           (dut_hip_status_rx_par_err),                             //                    .rx_par_err
		.tx_par_err           (dut_hip_status_tx_par_err),                             //                    .tx_par_err
		.cfg_par_err          (dut_hip_status_cfg_par_err),                            //                    .cfg_par_err
		.ko_cpl_spc_header    (dut_hip_status_ko_cpl_spc_header),                      //                    .ko_cpl_spc_header
		.ko_cpl_spc_data      (dut_hip_status_ko_cpl_spc_data),                        //                    .ko_cpl_spc_data
		.currentspeed         (dut_hip_currentspeed_currentspeed),                     //    hip_currentspeed.currentspeed
		.reconfig_to_xcvr     (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (dut_reconfig_from_xcvr_reconfig_from_xcvr),             //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (),                                                      // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (hip_serial_rx_in0),                                     //          hip_serial.rx_in0
		.rx_in1               (hip_serial_rx_in1),                                     //                    .rx_in1
		.rx_in2               (hip_serial_rx_in2),                                     //                    .rx_in2
		.rx_in3               (hip_serial_rx_in3),                                     //                    .rx_in3
		.tx_out0              (hip_serial_tx_out0),                                    //                    .tx_out0
		.tx_out1              (hip_serial_tx_out1),                                    //                    .tx_out1
		.tx_out2              (hip_serial_tx_out2),                                    //                    .tx_out2
		.tx_out3              (hip_serial_tx_out3),                                    //                    .tx_out3
		.sim_pipe_pclk_in     (),                                                      //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (),                                                      //                    .sim_pipe_rate
		.sim_ltssmstate       (),                                                      //                    .sim_ltssmstate
		.eidleinfersel0       (),                                                      //                    .eidleinfersel0
		.eidleinfersel1       (),                                                      //                    .eidleinfersel1
		.eidleinfersel2       (),                                                      //                    .eidleinfersel2
		.eidleinfersel3       (),                                                      //                    .eidleinfersel3
		.powerdown0           (),                                                      //                    .powerdown0
		.powerdown1           (),                                                      //                    .powerdown1
		.powerdown2           (),                                                      //                    .powerdown2
		.powerdown3           (),                                                      //                    .powerdown3
		.rxpolarity0          (),                                                      //                    .rxpolarity0
		.rxpolarity1          (),                                                      //                    .rxpolarity1
		.rxpolarity2          (),                                                      //                    .rxpolarity2
		.rxpolarity3          (),                                                      //                    .rxpolarity3
		.txcompl0             (),                                                      //                    .txcompl0
		.txcompl1             (),                                                      //                    .txcompl1
		.txcompl2             (),                                                      //                    .txcompl2
		.txcompl3             (),                                                      //                    .txcompl3
		.txdata0              (),                                                      //                    .txdata0
		.txdata1              (),                                                      //                    .txdata1
		.txdata2              (),                                                      //                    .txdata2
		.txdata3              (),                                                      //                    .txdata3
		.txdatak0             (),                                                      //                    .txdatak0
		.txdatak1             (),                                                      //                    .txdatak1
		.txdatak2             (),                                                      //                    .txdatak2
		.txdatak3             (),                                                      //                    .txdatak3
		.txdetectrx0          (),                                                      //                    .txdetectrx0
		.txdetectrx1          (),                                                      //                    .txdetectrx1
		.txdetectrx2          (),                                                      //                    .txdetectrx2
		.txdetectrx3          (),                                                      //                    .txdetectrx3
		.txelecidle0          (),                                                      //                    .txelecidle0
		.txelecidle1          (),                                                      //                    .txelecidle1
		.txelecidle2          (),                                                      //                    .txelecidle2
		.txelecidle3          (),                                                      //                    .txelecidle3
		.txdeemph0            (),                                                      //                    .txdeemph0
		.txdeemph1            (),                                                      //                    .txdeemph1
		.txdeemph2            (),                                                      //                    .txdeemph2
		.txdeemph3            (),                                                      //                    .txdeemph3
		.txmargin0            (),                                                      //                    .txmargin0
		.txmargin1            (),                                                      //                    .txmargin1
		.txmargin2            (),                                                      //                    .txmargin2
		.txmargin3            (),                                                      //                    .txmargin3
		.txswing0             (),                                                      //                    .txswing0
		.txswing1             (),                                                      //                    .txswing1
		.txswing2             (),                                                      //                    .txswing2
		.txswing3             (),                                                      //                    .txswing3
		.phystatus0           (),                                                      //                    .phystatus0
		.phystatus1           (),                                                      //                    .phystatus1
		.phystatus2           (),                                                      //                    .phystatus2
		.phystatus3           (),                                                      //                    .phystatus3
		.rxdata0              (),                                                      //                    .rxdata0
		.rxdata1              (),                                                      //                    .rxdata1
		.rxdata2              (),                                                      //                    .rxdata2
		.rxdata3              (),                                                      //                    .rxdata3
		.rxdatak0             (),                                                      //                    .rxdatak0
		.rxdatak1             (),                                                      //                    .rxdatak1
		.rxdatak2             (),                                                      //                    .rxdatak2
		.rxdatak3             (),                                                      //                    .rxdatak3
		.rxelecidle0          (),                                                      //                    .rxelecidle0
		.rxelecidle1          (),                                                      //                    .rxelecidle1
		.rxelecidle2          (),                                                      //                    .rxelecidle2
		.rxelecidle3          (),                                                      //                    .rxelecidle3
		.rxstatus0            (),                                                      //                    .rxstatus0
		.rxstatus1            (),                                                      //                    .rxstatus1
		.rxstatus2            (),                                                      //                    .rxstatus2
		.rxstatus3            (),                                                      //                    .rxstatus3
		.rxvalid0             (),                                                      //                    .rxvalid0
		.rxvalid1             (),                                                      //                    .rxvalid1
		.rxvalid2             (),                                                      //                    .rxvalid2
		.rxvalid3             (),                                                      //                    .rxvalid3
		.test_in              (hip_ctrl_test_in),                                      //            hip_ctrl.test_in
		.simu_mode_pipe       (hip_ctrl_simu_mode_pipe),                               //                    .simu_mode_pipe
		.TxsChipSelect_i      (),                                                      //                 Txs.chipselect
		.TxsByteEnable_i      (),                                                      //                    .byteenable
		.TxsReadData_o        (),                                                      //                    .readdata
		.TxsWriteData_i       (),                                                      //                    .writedata
		.TxsRead_i            (),                                                      //                    .read
		.TxsWrite_i           (),                                                      //                    .write
		.TxsBurstCount_i      (),                                                      //                    .burstcount
		.TxsReadDataValid_o   (),                                                      //                    .readdatavalid
		.TxsWaitRequest_o     (),                                                      //                    .waitrequest
		.TxsAddress_i         (),                                                      //                    .address
		.CraChipSelect_i      (mm_interconnect_0_dut_cra_chipselect),                  //                 Cra.chipselect
		.CraAddress_i         (mm_interconnect_0_dut_cra_address),                     //                    .address
		.CraByteEnable_i      (mm_interconnect_0_dut_cra_byteenable),                  //                    .byteenable
		.CraRead              (mm_interconnect_0_dut_cra_read),                        //                    .read
		.CraReadData_o        (mm_interconnect_0_dut_cra_readdata),                    //                    .readdata
		.CraWrite             (mm_interconnect_0_dut_cra_write),                       //                    .write
		.CraWriteData_i       (mm_interconnect_0_dut_cra_writedata),                   //                    .writedata
		.CraWaitRequest_o     (mm_interconnect_0_dut_cra_waitrequest),                 //                    .waitrequest
		.CraIrq_o             (),                                                      //              CraIrq.irq
		.rx_in4               (1'b0),                                                  //         (terminated)
		.rx_in5               (1'b0),                                                  //         (terminated)
		.rx_in6               (1'b0),                                                  //         (terminated)
		.rx_in7               (1'b0),                                                  //         (terminated)
		.tx_out4              (),                                                      //         (terminated)
		.tx_out5              (),                                                      //         (terminated)
		.tx_out6              (),                                                      //         (terminated)
		.tx_out7              (),                                                      //         (terminated)
		.eidleinfersel4       (),                                                      //         (terminated)
		.eidleinfersel5       (),                                                      //         (terminated)
		.eidleinfersel6       (),                                                      //         (terminated)
		.eidleinfersel7       (),                                                      //         (terminated)
		.powerdown4           (),                                                      //         (terminated)
		.powerdown5           (),                                                      //         (terminated)
		.powerdown6           (),                                                      //         (terminated)
		.powerdown7           (),                                                      //         (terminated)
		.rxpolarity4          (),                                                      //         (terminated)
		.rxpolarity5          (),                                                      //         (terminated)
		.rxpolarity6          (),                                                      //         (terminated)
		.rxpolarity7          (),                                                      //         (terminated)
		.txcompl4             (),                                                      //         (terminated)
		.txcompl5             (),                                                      //         (terminated)
		.txcompl6             (),                                                      //         (terminated)
		.txcompl7             (),                                                      //         (terminated)
		.txdata4              (),                                                      //         (terminated)
		.txdata5              (),                                                      //         (terminated)
		.txdata6              (),                                                      //         (terminated)
		.txdata7              (),                                                      //         (terminated)
		.txdatak4             (),                                                      //         (terminated)
		.txdatak5             (),                                                      //         (terminated)
		.txdatak6             (),                                                      //         (terminated)
		.txdatak7             (),                                                      //         (terminated)
		.txdetectrx4          (),                                                      //         (terminated)
		.txdetectrx5          (),                                                      //         (terminated)
		.txdetectrx6          (),                                                      //         (terminated)
		.txdetectrx7          (),                                                      //         (terminated)
		.txelecidle4          (),                                                      //         (terminated)
		.txelecidle5          (),                                                      //         (terminated)
		.txelecidle6          (),                                                      //         (terminated)
		.txelecidle7          (),                                                      //         (terminated)
		.txdeemph4            (),                                                      //         (terminated)
		.txdeemph5            (),                                                      //         (terminated)
		.txdeemph6            (),                                                      //         (terminated)
		.txdeemph7            (),                                                      //         (terminated)
		.txmargin4            (),                                                      //         (terminated)
		.txmargin5            (),                                                      //         (terminated)
		.txmargin6            (),                                                      //         (terminated)
		.txmargin7            (),                                                      //         (terminated)
		.txswing4             (),                                                      //         (terminated)
		.txswing5             (),                                                      //         (terminated)
		.txswing6             (),                                                      //         (terminated)
		.txswing7             (),                                                      //         (terminated)
		.phystatus4           (1'b0),                                                  //         (terminated)
		.phystatus5           (1'b0),                                                  //         (terminated)
		.phystatus6           (1'b0),                                                  //         (terminated)
		.phystatus7           (1'b0),                                                  //         (terminated)
		.rxdata4              (8'b00000000),                                           //         (terminated)
		.rxdata5              (8'b00000000),                                           //         (terminated)
		.rxdata6              (8'b00000000),                                           //         (terminated)
		.rxdata7              (8'b00000000),                                           //         (terminated)
		.rxdatak4             (1'b0),                                                  //         (terminated)
		.rxdatak5             (1'b0),                                                  //         (terminated)
		.rxdatak6             (1'b0),                                                  //         (terminated)
		.rxdatak7             (1'b0),                                                  //         (terminated)
		.rxelecidle4          (1'b0),                                                  //         (terminated)
		.rxelecidle5          (1'b0),                                                  //         (terminated)
		.rxelecidle6          (1'b0),                                                  //         (terminated)
		.rxelecidle7          (1'b0),                                                  //         (terminated)
		.rxstatus4            (3'b000),                                                //         (terminated)
		.rxstatus5            (3'b000),                                                //         (terminated)
		.rxstatus6            (3'b000),                                                //         (terminated)
		.rxstatus7            (3'b000),                                                //         (terminated)
		.rxvalid4             (1'b0),                                                  //         (terminated)
		.rxvalid5             (1'b0),                                                  //         (terminated)
		.rxvalid6             (1'b0),                                                  //         (terminated)
		.rxvalid7             (1'b0),                                                  //         (terminated)
		.rxdataskip0          (1'b0),                                                  //         (terminated)
		.rxdataskip1          (1'b0),                                                  //         (terminated)
		.rxdataskip2          (1'b0),                                                  //         (terminated)
		.rxdataskip3          (1'b0),                                                  //         (terminated)
		.rxdataskip4          (1'b0),                                                  //         (terminated)
		.rxdataskip5          (1'b0),                                                  //         (terminated)
		.rxdataskip6          (1'b0),                                                  //         (terminated)
		.rxdataskip7          (1'b0),                                                  //         (terminated)
		.rxblkst0             (1'b0),                                                  //         (terminated)
		.rxblkst1             (1'b0),                                                  //         (terminated)
		.rxblkst2             (1'b0),                                                  //         (terminated)
		.rxblkst3             (1'b0),                                                  //         (terminated)
		.rxblkst4             (1'b0),                                                  //         (terminated)
		.rxblkst5             (1'b0),                                                  //         (terminated)
		.rxblkst6             (1'b0),                                                  //         (terminated)
		.rxblkst7             (1'b0),                                                  //         (terminated)
		.rxsynchd0            (2'b00),                                                 //         (terminated)
		.rxsynchd1            (2'b00),                                                 //         (terminated)
		.rxsynchd2            (2'b00),                                                 //         (terminated)
		.rxsynchd3            (2'b00),                                                 //         (terminated)
		.rxsynchd4            (2'b00),                                                 //         (terminated)
		.rxsynchd5            (2'b00),                                                 //         (terminated)
		.rxsynchd6            (2'b00),                                                 //         (terminated)
		.rxsynchd7            (2'b00),                                                 //         (terminated)
		.rxfreqlocked0        (1'b0),                                                  //         (terminated)
		.rxfreqlocked1        (1'b0),                                                  //         (terminated)
		.rxfreqlocked2        (1'b0),                                                  //         (terminated)
		.rxfreqlocked3        (1'b0),                                                  //         (terminated)
		.rxfreqlocked4        (1'b0),                                                  //         (terminated)
		.rxfreqlocked5        (1'b0),                                                  //         (terminated)
		.rxfreqlocked6        (1'b0),                                                  //         (terminated)
		.rxfreqlocked7        (1'b0),                                                  //         (terminated)
		.currentcoeff0        (),                                                      //         (terminated)
		.currentcoeff1        (),                                                      //         (terminated)
		.currentcoeff2        (),                                                      //         (terminated)
		.currentcoeff3        (),                                                      //         (terminated)
		.currentcoeff4        (),                                                      //         (terminated)
		.currentcoeff5        (),                                                      //         (terminated)
		.currentcoeff6        (),                                                      //         (terminated)
		.currentcoeff7        (),                                                      //         (terminated)
		.currentrxpreset0     (),                                                      //         (terminated)
		.currentrxpreset1     (),                                                      //         (terminated)
		.currentrxpreset2     (),                                                      //         (terminated)
		.currentrxpreset3     (),                                                      //         (terminated)
		.currentrxpreset4     (),                                                      //         (terminated)
		.currentrxpreset5     (),                                                      //         (terminated)
		.currentrxpreset6     (),                                                      //         (terminated)
		.currentrxpreset7     (),                                                      //         (terminated)
		.txsynchd0            (),                                                      //         (terminated)
		.txsynchd1            (),                                                      //         (terminated)
		.txsynchd2            (),                                                      //         (terminated)
		.txsynchd3            (),                                                      //         (terminated)
		.txsynchd4            (),                                                      //         (terminated)
		.txsynchd5            (),                                                      //         (terminated)
		.txsynchd6            (),                                                      //         (terminated)
		.txsynchd7            (),                                                      //         (terminated)
		.txblkst0             (),                                                      //         (terminated)
		.txblkst1             (),                                                      //         (terminated)
		.txblkst2             (),                                                      //         (terminated)
		.txblkst3             (),                                                      //         (terminated)
		.txblkst4             (),                                                      //         (terminated)
		.txblkst5             (),                                                      //         (terminated)
		.txblkst6             (),                                                      //         (terminated)
		.txblkst7             ()                                                       //         (terminated)
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (6),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (1),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),       //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (mgmt_clk_clk),                                          //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (mgmt_rst_reset),                                        //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),          //      reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),             //                   .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),         //                   .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest),      //                   .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),            //                   .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),        //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (dut_reconfig_from_xcvr_reconfig_from_xcvr),             // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                      //        (terminated)
		.rx_cal_busy               (),                                                      //        (terminated)
		.cal_busy_in               (1'b0),                                                  //        (terminated)
		.reconfig_mif_address      (),                                                      //        (terminated)
		.reconfig_mif_read         (),                                                      //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                  //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                   //        (terminated)
	);

	avl_to_asmi avl_to_asmi_0 (
		.avs_s0_address         (mm_interconnect_0_avl_to_asmi_0_s0_address),   //          s0.address
		.avs_s0_read            (mm_interconnect_0_avl_to_asmi_0_s0_read),      //            .read
		.avs_s0_readdata        (mm_interconnect_0_avl_to_asmi_0_s0_readdata),  //            .readdata
		.avs_s0_write           (mm_interconnect_0_avl_to_asmi_0_s0_write),     //            .write
		.avs_s0_writedata       (mm_interconnect_0_avl_to_asmi_0_s0_writedata), //            .writedata
		.clk                    (dut_coreclkout_clk),                           //       clock.clk
		.reset                  (rst_controller_reset_out_reset),               //       reset.reset
		.asmi_sfl_address       (avl_to_asmi_0_conduit_end_sfl_address),        // conduit_end.sfl_address
		.asmi_sfl_read          (avl_to_asmi_0_conduit_end_sfl_read),           //            .sfl_read
		.asmi_sfl_readdata_from (avl_to_asmi_0_conduit_end_sfl_readdata_from),  //            .sfl_readdata_from
		.asmi_sfl_write         (avl_to_asmi_0_conduit_end_sfl_write),          //            .sfl_write
		.asmi_sfl_writedata_to  (avl_to_asmi_0_conduit_end_sfl_writedata_to),   //            .sfl_writedata_to
		.asmi_sfl_clk           (avl_to_asmi_0_conduit_end_sfl_clk),            //            .sfl_clk
		.asmi_sfl_reset         (avl_to_asmi_0_conduit_end_sfl_reset)           //            .sfl_reset
	);

	pcie_hip_avmm_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk               (clk_clk),                                                     //      pll_ref_clk.clk
		.global_reset_n            (reset_reset_n),                                               //     global_reset.reset_n
		.soft_reset_n              (reset_reset_n),                                               //       soft_reset.reset_n
		.afi_clk                   (mem_if_ddr3_emif_0_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                                            //     afi_half_clk.clk
		.afi_reset_n               (),                                                            //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                            // afi_reset_export.reset_n
		.mem_a                     (memory_mem_a),                                                //           memory.mem_a
		.mem_ba                    (memory_mem_ba),                                               //                 .mem_ba
		.mem_ck                    (memory_mem_ck),                                               //                 .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                                             //                 .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                              //                 .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                                             //                 .mem_cs_n
		.mem_dm                    (memory_mem_dm),                                               //                 .mem_dm
		.mem_ras_n                 (memory_mem_ras_n),                                            //                 .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                                            //                 .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                                             //                 .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                                          //                 .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                               //                 .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                              //                 .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                                            //                 .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                              //                 .mem_odt
		.avl_ready                 (mm_interconnect_1_mem_if_ddr3_emif_0_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_1_mem_if_ddr3_emif_0_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_1_mem_if_ddr3_emif_0_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_1_mem_if_ddr3_emif_0_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_1_mem_if_ddr3_emif_0_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_1_mem_if_ddr3_emif_0_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_1_mem_if_ddr3_emif_0_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_1_mem_if_ddr3_emif_0_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_1_mem_if_ddr3_emif_0_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_1_mem_if_ddr3_emif_0_avl_burstcount),         //                 .burstcount
		.local_init_done           (),                                                            //           status.local_init_done
		.local_cal_success         (),                                                            //                 .local_cal_success
		.local_cal_fail            (),                                                            //                 .local_cal_fail
		.oct_rzqin                 (oct_rzqin),                                                   //              oct.rzqin
		.pll_mem_clk               (),                                                            //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                                            //                 .pll_write_clk
		.pll_locked                (),                                                            //                 .pll_locked
		.pll_write_clk_pre_phy_clk (),                                                            //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                                            //                 .pll_addr_cmd_clk
		.pll_avl_clk               (),                                                            //                 .pll_avl_clk
		.pll_config_clk            (),                                                            //                 .pll_config_clk
		.pll_hr_clk                (),                                                            //                 .pll_hr_clk
		.pll_p2c_read_clk          (),                                                            //                 .pll_p2c_read_clk
		.pll_c2p_write_clk         (),                                                            //                 .pll_c2p_write_clk
		.csr_addr                  (mm_interconnect_0_mem_if_ddr3_emif_0_csr_address),            //              csr.address
		.csr_read_req              (mm_interconnect_0_mem_if_ddr3_emif_0_csr_read),               //                 .read
		.csr_rdata                 (mm_interconnect_0_mem_if_ddr3_emif_0_csr_readdata),           //                 .readdata
		.csr_write_req             (mm_interconnect_0_mem_if_ddr3_emif_0_csr_write),              //                 .write
		.csr_wdata                 (mm_interconnect_0_mem_if_ddr3_emif_0_csr_writedata),          //                 .writedata
		.csr_waitrequest           (mm_interconnect_0_mem_if_ddr3_emif_0_csr_waitrequest),        //                 .waitrequest
		.csr_be                    (mm_interconnect_0_mem_if_ddr3_emif_0_csr_byteenable),         //                 .byteenable
		.csr_rdata_valid           (mm_interconnect_0_mem_if_ddr3_emif_0_csr_readdatavalid),      //                 .readdatavalid
		.seq_debug_addr            (),                                                            //        seq_debug.address
		.seq_debug_read_req        (),                                                            //                 .read
		.seq_debug_rdata           (),                                                            //                 .readdata
		.seq_debug_write_req       (),                                                            //                 .write
		.seq_debug_wdata           (),                                                            //                 .writedata
		.seq_debug_waitrequest     (),                                                            //                 .waitrequest
		.seq_debug_be              (),                                                            //                 .byteenable
		.seq_debug_rdata_valid     ()                                                             //                 .readdatavalid
	);

	pcie_hip_avmm_mem_if_ddr3_emif_0 mem_if_ddr3_emif_1 (
		.pll_ref_clk               (clk_1_clk),                                                   //      pll_ref_clk.clk
		.global_reset_n            (reset_1_reset_n),                                             //     global_reset.reset_n
		.soft_reset_n              (reset_1_reset_n),                                             //       soft_reset.reset_n
		.afi_clk                   (mem_if_ddr3_emif_1_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                                            //     afi_half_clk.clk
		.afi_reset_n               (),                                                            //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                            // afi_reset_export.reset_n
		.mem_a                     (memory_1_mem_a),                                              //           memory.mem_a
		.mem_ba                    (memory_1_mem_ba),                                             //                 .mem_ba
		.mem_ck                    (memory_1_mem_ck),                                             //                 .mem_ck
		.mem_ck_n                  (memory_1_mem_ck_n),                                           //                 .mem_ck_n
		.mem_cke                   (memory_1_mem_cke),                                            //                 .mem_cke
		.mem_cs_n                  (memory_1_mem_cs_n),                                           //                 .mem_cs_n
		.mem_dm                    (memory_1_mem_dm),                                             //                 .mem_dm
		.mem_ras_n                 (memory_1_mem_ras_n),                                          //                 .mem_ras_n
		.mem_cas_n                 (memory_1_mem_cas_n),                                          //                 .mem_cas_n
		.mem_we_n                  (memory_1_mem_we_n),                                           //                 .mem_we_n
		.mem_reset_n               (memory_1_mem_reset_n),                                        //                 .mem_reset_n
		.mem_dq                    (memory_1_mem_dq),                                             //                 .mem_dq
		.mem_dqs                   (memory_1_mem_dqs),                                            //                 .mem_dqs
		.mem_dqs_n                 (memory_1_mem_dqs_n),                                          //                 .mem_dqs_n
		.mem_odt                   (memory_1_mem_odt),                                            //                 .mem_odt
		.avl_ready                 (mm_interconnect_2_mem_if_ddr3_emif_1_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_2_mem_if_ddr3_emif_1_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_2_mem_if_ddr3_emif_1_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_2_mem_if_ddr3_emif_1_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_2_mem_if_ddr3_emif_1_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_2_mem_if_ddr3_emif_1_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_2_mem_if_ddr3_emif_1_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_2_mem_if_ddr3_emif_1_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_2_mem_if_ddr3_emif_1_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_2_mem_if_ddr3_emif_1_avl_burstcount),         //                 .burstcount
		.local_init_done           (),                                                            //           status.local_init_done
		.local_cal_success         (),                                                            //                 .local_cal_success
		.local_cal_fail            (),                                                            //                 .local_cal_fail
		.oct_rzqin                 (oct_1_rzqin),                                                 //              oct.rzqin
		.pll_mem_clk               (),                                                            //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                                            //                 .pll_write_clk
		.pll_locked                (),                                                            //                 .pll_locked
		.pll_write_clk_pre_phy_clk (),                                                            //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                                            //                 .pll_addr_cmd_clk
		.pll_avl_clk               (),                                                            //                 .pll_avl_clk
		.pll_config_clk            (),                                                            //                 .pll_config_clk
		.pll_hr_clk                (),                                                            //                 .pll_hr_clk
		.pll_p2c_read_clk          (),                                                            //                 .pll_p2c_read_clk
		.pll_c2p_write_clk         (),                                                            //                 .pll_c2p_write_clk
		.csr_addr                  (mm_interconnect_0_mem_if_ddr3_emif_1_csr_address),            //              csr.address
		.csr_read_req              (mm_interconnect_0_mem_if_ddr3_emif_1_csr_read),               //                 .read
		.csr_rdata                 (mm_interconnect_0_mem_if_ddr3_emif_1_csr_readdata),           //                 .readdata
		.csr_write_req             (mm_interconnect_0_mem_if_ddr3_emif_1_csr_write),              //                 .write
		.csr_wdata                 (mm_interconnect_0_mem_if_ddr3_emif_1_csr_writedata),          //                 .writedata
		.csr_waitrequest           (mm_interconnect_0_mem_if_ddr3_emif_1_csr_waitrequest),        //                 .waitrequest
		.csr_be                    (mm_interconnect_0_mem_if_ddr3_emif_1_csr_byteenable),         //                 .byteenable
		.csr_rdata_valid           (mm_interconnect_0_mem_if_ddr3_emif_1_csr_readdatavalid),      //                 .readdatavalid
		.seq_debug_addr            (),                                                            //        seq_debug.address
		.seq_debug_read_req        (),                                                            //                 .read
		.seq_debug_rdata           (),                                                            //                 .readdata
		.seq_debug_write_req       (),                                                            //                 .write
		.seq_debug_wdata           (),                                                            //                 .writedata
		.seq_debug_waitrequest     (),                                                            //                 .waitrequest
		.seq_debug_be              (),                                                            //                 .byteenable
		.seq_debug_rdata_valid     ()                                                             //                 .readdatavalid
	);

	altpcie_reconfig_driver #(
		.INTENDED_DEVICE_FAMILY        ("Stratix V"),
		.gen123_lane_rate_mode_hwtcl   ("Gen3 (8.0 Gbps)"),
		.number_of_reconfig_interfaces (6)
	) pcie_reconfig_driver_0 (
		.reconfig_xcvr_clk         (reconfig_xcvr_clk_clk),                            // reconfig_xcvr_clk.clk
		.reconfig_xcvr_rst         (reconfig_xcvr_rst_reset),                          // reconfig_xcvr_rst.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),     //     reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),        //                  .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),    //                  .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest), //                  .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),       //                  .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),   //                  .writedata
		.currentspeed              (dut_hip_currentspeed_currentspeed),                //  hip_currentspeed.currentspeed
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),  //     reconfig_busy.reconfig_busy
		.pld_clk                   (dut_coreclkout_clk),                               //           pld_clk.clk
		.derr_cor_ext_rcv_drv      (dut_hip_status_derr_cor_ext_rcv),                  //    hip_status_drv.derr_cor_ext_rcv
		.derr_cor_ext_rpl_drv      (dut_hip_status_derr_cor_ext_rpl),                  //                  .derr_cor_ext_rpl
		.derr_rpl_drv              (dut_hip_status_derr_rpl),                          //                  .derr_rpl
		.dlup_exit_drv             (dut_hip_status_dlup_exit),                         //                  .dlup_exit
		.ev128ns_drv               (dut_hip_status_ev128ns),                           //                  .ev128ns
		.ev1us_drv                 (dut_hip_status_ev1us),                             //                  .ev1us
		.hotrst_exit_drv           (dut_hip_status_hotrst_exit),                       //                  .hotrst_exit
		.int_status_drv            (dut_hip_status_int_status),                        //                  .int_status
		.l2_exit_drv               (dut_hip_status_l2_exit),                           //                  .l2_exit
		.lane_act_drv              (dut_hip_status_lane_act),                          //                  .lane_act
		.ltssmstate_drv            (dut_hip_status_ltssmstate),                        //                  .ltssmstate
		.dlup_drv                  (dut_hip_status_dlup),                              //                  .dlup
		.rx_par_err_drv            (dut_hip_status_rx_par_err),                        //                  .rx_par_err
		.tx_par_err_drv            (dut_hip_status_tx_par_err),                        //                  .tx_par_err
		.cfg_par_err_drv           (dut_hip_status_cfg_par_err),                       //                  .cfg_par_err
		.ko_cpl_spc_header_drv     (dut_hip_status_ko_cpl_spc_header),                 //                  .ko_cpl_spc_header
		.ko_cpl_spc_data_drv       (dut_hip_status_ko_cpl_spc_data),                   //                  .ko_cpl_spc_data
		.cal_busy_in               ()                                                  //       (terminated)
	);

	pcie_hip_avmm_mm_interconnect_0 mm_interconnect_0 (
		.DUT_coreclkout_clk                                                  (dut_coreclkout_clk),                                     //                                                DUT_coreclkout.clk
		.mem_if_ddr3_emif_0_afi_clk_clk                                      (mem_if_ddr3_emif_0_afi_clk_clk),                         //                                    mem_if_ddr3_emif_0_afi_clk.clk
		.mem_if_ddr3_emif_1_afi_clk_clk                                      (mem_if_ddr3_emif_1_afi_clk_clk),                         //                                    mem_if_ddr3_emif_1_afi_clk.clk
		.avl_to_asmi_0_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                         //                     avl_to_asmi_0_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_csr_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                     // mem_if_ddr3_emif_0_csr_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                     //           mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_1_csr_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                     // mem_if_ddr3_emif_1_csr_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_1_soft_reset_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                     //           mem_if_ddr3_emif_1_soft_reset_reset_bridge_in_reset.reset
		.DUT_Rxm_BAR0_address                                                (dut_rxm_bar0_address),                                   //                                                  DUT_Rxm_BAR0.address
		.DUT_Rxm_BAR0_waitrequest                                            (dut_rxm_bar0_waitrequest),                               //                                                              .waitrequest
		.DUT_Rxm_BAR0_burstcount                                             (dut_rxm_bar0_burstcount),                                //                                                              .burstcount
		.DUT_Rxm_BAR0_byteenable                                             (dut_rxm_bar0_byteenable),                                //                                                              .byteenable
		.DUT_Rxm_BAR0_read                                                   (dut_rxm_bar0_read),                                      //                                                              .read
		.DUT_Rxm_BAR0_readdata                                               (dut_rxm_bar0_readdata),                                  //                                                              .readdata
		.DUT_Rxm_BAR0_readdatavalid                                          (dut_rxm_bar0_readdatavalid),                             //                                                              .readdatavalid
		.DUT_Rxm_BAR0_write                                                  (dut_rxm_bar0_write),                                     //                                                              .write
		.DUT_Rxm_BAR0_writedata                                              (dut_rxm_bar0_writedata),                                 //                                                              .writedata
		.avl_to_asmi_0_s0_address                                            (mm_interconnect_0_avl_to_asmi_0_s0_address),             //                                              avl_to_asmi_0_s0.address
		.avl_to_asmi_0_s0_write                                              (mm_interconnect_0_avl_to_asmi_0_s0_write),               //                                                              .write
		.avl_to_asmi_0_s0_read                                               (mm_interconnect_0_avl_to_asmi_0_s0_read),                //                                                              .read
		.avl_to_asmi_0_s0_readdata                                           (mm_interconnect_0_avl_to_asmi_0_s0_readdata),            //                                                              .readdata
		.avl_to_asmi_0_s0_writedata                                          (mm_interconnect_0_avl_to_asmi_0_s0_writedata),           //                                                              .writedata
		.DUT_Cra_address                                                     (mm_interconnect_0_dut_cra_address),                      //                                                       DUT_Cra.address
		.DUT_Cra_write                                                       (mm_interconnect_0_dut_cra_write),                        //                                                              .write
		.DUT_Cra_read                                                        (mm_interconnect_0_dut_cra_read),                         //                                                              .read
		.DUT_Cra_readdata                                                    (mm_interconnect_0_dut_cra_readdata),                     //                                                              .readdata
		.DUT_Cra_writedata                                                   (mm_interconnect_0_dut_cra_writedata),                    //                                                              .writedata
		.DUT_Cra_byteenable                                                  (mm_interconnect_0_dut_cra_byteenable),                   //                                                              .byteenable
		.DUT_Cra_waitrequest                                                 (mm_interconnect_0_dut_cra_waitrequest),                  //                                                              .waitrequest
		.DUT_Cra_chipselect                                                  (mm_interconnect_0_dut_cra_chipselect),                   //                                                              .chipselect
		.mem_if_ddr3_emif_0_csr_address                                      (mm_interconnect_0_mem_if_ddr3_emif_0_csr_address),       //                                        mem_if_ddr3_emif_0_csr.address
		.mem_if_ddr3_emif_0_csr_write                                        (mm_interconnect_0_mem_if_ddr3_emif_0_csr_write),         //                                                              .write
		.mem_if_ddr3_emif_0_csr_read                                         (mm_interconnect_0_mem_if_ddr3_emif_0_csr_read),          //                                                              .read
		.mem_if_ddr3_emif_0_csr_readdata                                     (mm_interconnect_0_mem_if_ddr3_emif_0_csr_readdata),      //                                                              .readdata
		.mem_if_ddr3_emif_0_csr_writedata                                    (mm_interconnect_0_mem_if_ddr3_emif_0_csr_writedata),     //                                                              .writedata
		.mem_if_ddr3_emif_0_csr_byteenable                                   (mm_interconnect_0_mem_if_ddr3_emif_0_csr_byteenable),    //                                                              .byteenable
		.mem_if_ddr3_emif_0_csr_readdatavalid                                (mm_interconnect_0_mem_if_ddr3_emif_0_csr_readdatavalid), //                                                              .readdatavalid
		.mem_if_ddr3_emif_0_csr_waitrequest                                  (mm_interconnect_0_mem_if_ddr3_emif_0_csr_waitrequest),   //                                                              .waitrequest
		.mem_if_ddr3_emif_1_csr_address                                      (mm_interconnect_0_mem_if_ddr3_emif_1_csr_address),       //                                        mem_if_ddr3_emif_1_csr.address
		.mem_if_ddr3_emif_1_csr_write                                        (mm_interconnect_0_mem_if_ddr3_emif_1_csr_write),         //                                                              .write
		.mem_if_ddr3_emif_1_csr_read                                         (mm_interconnect_0_mem_if_ddr3_emif_1_csr_read),          //                                                              .read
		.mem_if_ddr3_emif_1_csr_readdata                                     (mm_interconnect_0_mem_if_ddr3_emif_1_csr_readdata),      //                                                              .readdata
		.mem_if_ddr3_emif_1_csr_writedata                                    (mm_interconnect_0_mem_if_ddr3_emif_1_csr_writedata),     //                                                              .writedata
		.mem_if_ddr3_emif_1_csr_byteenable                                   (mm_interconnect_0_mem_if_ddr3_emif_1_csr_byteenable),    //                                                              .byteenable
		.mem_if_ddr3_emif_1_csr_readdatavalid                                (mm_interconnect_0_mem_if_ddr3_emif_1_csr_readdatavalid), //                                                              .readdatavalid
		.mem_if_ddr3_emif_1_csr_waitrequest                                  (mm_interconnect_0_mem_if_ddr3_emif_1_csr_waitrequest)    //                                                              .waitrequest
	);

	pcie_hip_avmm_mm_interconnect_1 mm_interconnect_1 (
		.DUT_coreclkout_clk                                                  (dut_coreclkout_clk),                                          //                                                DUT_coreclkout.clk
		.mem_if_ddr3_emif_0_afi_clk_clk                                      (mem_if_ddr3_emif_0_afi_clk_clk),                              //                                    mem_if_ddr3_emif_0_afi_clk.clk
		.mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                          //           mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset.reset
		.move_engine_0_rst_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                              //                       move_engine_0_rst_reset_bridge_in_reset.reset
		.DUT_Rxm_BAR2_address                                                (dut_rxm_bar2_address),                                        //                                                  DUT_Rxm_BAR2.address
		.DUT_Rxm_BAR2_waitrequest                                            (dut_rxm_bar2_waitrequest),                                    //                                                              .waitrequest
		.DUT_Rxm_BAR2_burstcount                                             (dut_rxm_bar2_burstcount),                                     //                                                              .burstcount
		.DUT_Rxm_BAR2_byteenable                                             (dut_rxm_bar2_byteenable),                                     //                                                              .byteenable
		.DUT_Rxm_BAR2_read                                                   (dut_rxm_bar2_read),                                           //                                                              .read
		.DUT_Rxm_BAR2_readdata                                               (dut_rxm_bar2_readdata),                                       //                                                              .readdata
		.DUT_Rxm_BAR2_readdatavalid                                          (dut_rxm_bar2_readdatavalid),                                  //                                                              .readdatavalid
		.DUT_Rxm_BAR2_write                                                  (dut_rxm_bar2_write),                                          //                                                              .write
		.DUT_Rxm_BAR2_writedata                                              (dut_rxm_bar2_writedata),                                      //                                                              .writedata
		.move_engine_0_fast_master_address                                   (fast_mem_address),                                            //                                     move_engine_0_fast_master.address
		.move_engine_0_fast_master_waitrequest                               (fast_mem_waitrequest),                                        //                                                              .waitrequest
		.move_engine_0_fast_master_burstcount                                (fast_mem_burstcount),                                         //                                                              .burstcount
		.move_engine_0_fast_master_read                                      (fast_mem_read),                                               //                                                              .read
		.move_engine_0_fast_master_readdata                                  (fast_mem_readdata),                                           //                                                              .readdata
		.move_engine_0_fast_master_readdatavalid                             (fast_mem_readdatavalid),                                      //                                                              .readdatavalid
		.move_engine_0_fast_master_write                                     (fast_mem_write),                                              //                                                              .write
		.move_engine_0_fast_master_writedata                                 (fast_mem_writedata),                                          //                                                              .writedata
		.move_engine_0_fast_master_lock                                      (fast_mem_lock),                                               //                                                              .lock
		.mem_if_ddr3_emif_0_avl_address                                      (mm_interconnect_1_mem_if_ddr3_emif_0_avl_address),            //                                        mem_if_ddr3_emif_0_avl.address
		.mem_if_ddr3_emif_0_avl_write                                        (mm_interconnect_1_mem_if_ddr3_emif_0_avl_write),              //                                                              .write
		.mem_if_ddr3_emif_0_avl_read                                         (mm_interconnect_1_mem_if_ddr3_emif_0_avl_read),               //                                                              .read
		.mem_if_ddr3_emif_0_avl_readdata                                     (mm_interconnect_1_mem_if_ddr3_emif_0_avl_readdata),           //                                                              .readdata
		.mem_if_ddr3_emif_0_avl_writedata                                    (mm_interconnect_1_mem_if_ddr3_emif_0_avl_writedata),          //                                                              .writedata
		.mem_if_ddr3_emif_0_avl_beginbursttransfer                           (mm_interconnect_1_mem_if_ddr3_emif_0_avl_beginbursttransfer), //                                                              .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_burstcount                                   (mm_interconnect_1_mem_if_ddr3_emif_0_avl_burstcount),         //                                                              .burstcount
		.mem_if_ddr3_emif_0_avl_byteenable                                   (mm_interconnect_1_mem_if_ddr3_emif_0_avl_byteenable),         //                                                              .byteenable
		.mem_if_ddr3_emif_0_avl_readdatavalid                                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_readdatavalid),      //                                                              .readdatavalid
		.mem_if_ddr3_emif_0_avl_waitrequest                                  (~mm_interconnect_1_mem_if_ddr3_emif_0_avl_waitrequest)        //                                                              .waitrequest
	);

	pcie_hip_avmm_mm_interconnect_2 mm_interconnect_2 (
		.DUT_coreclkout_clk                                                  (dut_coreclkout_clk),                                          //                                                DUT_coreclkout.clk
		.mem_if_ddr3_emif_1_afi_clk_clk                                      (mem_if_ddr3_emif_1_afi_clk_clk),                              //                                    mem_if_ddr3_emif_1_afi_clk.clk
		.mem_if_ddr3_emif_1_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // mem_if_ddr3_emif_1_avl_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_1_soft_reset_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                          //           mem_if_ddr3_emif_1_soft_reset_reset_bridge_in_reset.reset
		.move_engine_0_rst_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                              //                       move_engine_0_rst_reset_bridge_in_reset.reset
		.DUT_Rxm_BAR4_address                                                (dut_rxm_bar4_address),                                        //                                                  DUT_Rxm_BAR4.address
		.DUT_Rxm_BAR4_waitrequest                                            (dut_rxm_bar4_waitrequest),                                    //                                                              .waitrequest
		.DUT_Rxm_BAR4_burstcount                                             (dut_rxm_bar4_burstcount),                                     //                                                              .burstcount
		.DUT_Rxm_BAR4_byteenable                                             (dut_rxm_bar4_byteenable),                                     //                                                              .byteenable
		.DUT_Rxm_BAR4_read                                                   (dut_rxm_bar4_read),                                           //                                                              .read
		.DUT_Rxm_BAR4_readdata                                               (dut_rxm_bar4_readdata),                                       //                                                              .readdata
		.DUT_Rxm_BAR4_readdatavalid                                          (dut_rxm_bar4_readdatavalid),                                  //                                                              .readdatavalid
		.DUT_Rxm_BAR4_write                                                  (dut_rxm_bar4_write),                                          //                                                              .write
		.DUT_Rxm_BAR4_writedata                                              (dut_rxm_bar4_writedata),                                      //                                                              .writedata
		.move_engine_0_slow_master_address                                   (slow_mem_address),                                            //                                     move_engine_0_slow_master.address
		.move_engine_0_slow_master_waitrequest                               (slow_mem_waitrequest),                                        //                                                              .waitrequest
		.move_engine_0_slow_master_burstcount                                (slow_mem_burstcount),                                         //                                                              .burstcount
		.move_engine_0_slow_master_read                                      (slow_mem_read),                                               //                                                              .read
		.move_engine_0_slow_master_readdata                                  (slow_mem_readdata),                                           //                                                              .readdata
		.move_engine_0_slow_master_readdatavalid                             (slow_mem_readdatavalid),                                      //                                                              .readdatavalid
		.move_engine_0_slow_master_write                                     (slow_mem_write),                                              //                                                              .write
		.move_engine_0_slow_master_writedata                                 (slow_mem_writedata),                                          //                                                              .writedata
		.move_engine_0_slow_master_lock                                      (slow_mem_lock),                                               //                                                              .lock
		.mem_if_ddr3_emif_1_avl_address                                      (mm_interconnect_2_mem_if_ddr3_emif_1_avl_address),            //                                        mem_if_ddr3_emif_1_avl.address
		.mem_if_ddr3_emif_1_avl_write                                        (mm_interconnect_2_mem_if_ddr3_emif_1_avl_write),              //                                                              .write
		.mem_if_ddr3_emif_1_avl_read                                         (mm_interconnect_2_mem_if_ddr3_emif_1_avl_read),               //                                                              .read
		.mem_if_ddr3_emif_1_avl_readdata                                     (mm_interconnect_2_mem_if_ddr3_emif_1_avl_readdata),           //                                                              .readdata
		.mem_if_ddr3_emif_1_avl_writedata                                    (mm_interconnect_2_mem_if_ddr3_emif_1_avl_writedata),          //                                                              .writedata
		.mem_if_ddr3_emif_1_avl_beginbursttransfer                           (mm_interconnect_2_mem_if_ddr3_emif_1_avl_beginbursttransfer), //                                                              .beginbursttransfer
		.mem_if_ddr3_emif_1_avl_burstcount                                   (mm_interconnect_2_mem_if_ddr3_emif_1_avl_burstcount),         //                                                              .burstcount
		.mem_if_ddr3_emif_1_avl_byteenable                                   (mm_interconnect_2_mem_if_ddr3_emif_1_avl_byteenable),         //                                                              .byteenable
		.mem_if_ddr3_emif_1_avl_readdatavalid                                (mm_interconnect_2_mem_if_ddr3_emif_1_avl_readdatavalid),      //                                                              .readdatavalid
		.mem_if_ddr3_emif_1_avl_waitrequest                                  (~mm_interconnect_2_mem_if_ddr3_emif_1_avl_waitrequest)        //                                                              .waitrequest
	);

	pcie_hip_avmm_irq_mapper irq_mapper (
		.clk        (dut_coreclkout_clk),             //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (dut_rxmirq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~dut_nreset_status_reset),       // reset_in0.reset
		.clk            (dut_coreclkout_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_1_reset_n),                   // reset_in0.reset
		.clk            (mem_if_ddr3_emif_1_afi_clk_clk),     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
